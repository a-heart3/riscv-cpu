`ifndef PIPELINE_VH
    `define PIPELINE_VH

    `define BRANCH_DATA 33
    `define FS_DATA     64
    `define ID_DATA     91
    `define EX_DATA     80
    `define EX_MEM_DATA 42
    `define MEM_DATA    74

`endif