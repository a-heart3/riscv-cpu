`ifndef PIPELINE_VH
    `define PIPELINE_VH

    `define BRANCH_DATA 33
    `define FS_DATA     64

`endif