`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 05/10/2025 10:03:08 PM
// Design Name: 
// Module Name: data_ram
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module data_ram(
    input  [31:0] data_sram_addr,
    input  [31:0] data_sram_wdata,
    input         data_sram_en,
    input         data_sram_we,
    input  [ 2:0] data_sram_mode,
    input         data_sram_us,
    output [31:0] rdata
);


endmodule
