`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 05/06/2025 07:35:46 PM
// Design Name: 
// Module Name: top_tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module top_tb();
reg         clk;
reg         reset;
reg  [ 4:0] wb_rd;
reg  [31:0] wb_wdata;
reg         wb_we;
reg         mem_wb_reg_allow_in;
wire        mem_to_wb_reg_valid;
wire [73:0] mem_data;

top top(
    .clk                (clk                 ),
    .reset              (reset               ),
    .wb_rd              (wb_rd               ),
    .wb_wdata           (wb_wdata            ),
    .wb_we              (wb_we               ),
    .mem_wb_reg_allow_in(mem_wb_reg_allow_in ),
    .mem_to_wb_reg_valid(mem_to_wb_reg_valid ),
    .mem_data           (mem_data            )
);

initial begin
    clk <= 1'b0;
    reset <= 1'b1;
    wb_rd <= 5'b00001;
    wb_wdata <= 32'd1;
    wb_we <= 1'b1;
    mem_wb_reg_allow_in <= 1'b0;
    #10;
    reset <= 1'b0;
    mem_wb_reg_allow_in = 1'b1;
    wb_rd <= 5'b00010;
    wb_wdata <= 32'd2;
    wb_we <= 1'b1;
    #10;
    wb_we <= 1'b0;
end

always begin
    #5;
    clk <= ~clk;
end

endmodule
